.param var=0.000309
