TDO - TUNNEL DIODE OSCILLATOR	
VIN	3	0	0.399567
R1	2	3	0.2
LS  2 	1 	1UH	 IC=0.001044 
CS  1 	0 	1000PF
G1 1 0 	POLY(1)	1 0 0.084039 0.6 -1.5 1 	
.IC V(1)=-0.104675
.TRAN 1NS 5NS UIC
.PRINT V(1) I(LS) I(Vin)
.OPT BRIEF numdgt=10
.END
