.param var=-0.000664
