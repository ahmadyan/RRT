.param var=0.000955
