.param var=0