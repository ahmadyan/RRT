.param var=-0.000296
