.param var=0.000544
