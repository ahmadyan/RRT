.param var=0.000808
